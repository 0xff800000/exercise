$date
  Fri Nov 17 16:58:59 2017
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$var reg 1 ! clk_tb $end
$var reg 1 " res_tb $end
$var reg 4 # out_tb[3:0] $end
$scope module duv $end
$var reg 1 $ clk_i $end
$var reg 1 % rst_i $end
$var reg 1 & max_o $end
$var reg 4 ' out_o[3:0] $end
$var reg 4 ( current_state[3:0] $end
$var reg 4 ) next_state[3:0] $end
$upscope $end
$enddefinitions $end
#0
1!
1"
b0000 #
1$
1%
0&
b0000 '
bUUUU (
b0000 )
#10000000
0!
0"
0$
0%
#20000000
1!
b0001 #
1$
b0001 '
b0001 )
#30000000
0!
0$
#40000000
1!
b0011 #
1$
b0011 '
b0011 )
#50000000
0!
0$
#60000000
1!
b0111 #
1$
b0111 '
b0111 )
#70000000
0!
0$
#80000000
1!
b1111 #
1$
b1111 '
b1111 )
#90000000
0!
0$
#100000000
1!
b1110 #
1$
b1110 '
b1110 )
#110000000
0!
0$
#120000000
1!
b1100 #
1$
b1100 '
b1100 )
#130000000
0!
0$
#140000000
1!
b1000 #
1$
1&
b1000 '
b1000 )
#150000000
0!
0$
1&
#160000000
1!
b0000 #
1$
0&
b0000 '
b0000 )
#170000000
